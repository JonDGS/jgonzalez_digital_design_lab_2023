//module decoColor(
//		input logic [2:0] code,
//		output logic [7:0] r,
//		output logic [7:0] g,
//		output logic [7:0] b
//		);
//		
//	case(code)
//		0: begin
//			r <= 8'h00;
//			g <= 8'h00;
//			b <= 8'h00;
//		end
//		1: begin
//			r <= 8'h00;
//			g <= 8'h00;
//			b <= 8'h00;
//		end
//		2: begin
//			r <= 8'h00;
//			g <= 8'h00;
//			b <= 8'h00;
//		end
//		3: begin
//			r <= 8'h00;
//			g <= 8'h00;
//			b <= 8'h00;
//		end
//		4: begin
//			r <= 8'h00;
//			g <= 8'h00;
//			b <= 8'h00;
//		end
//		5: begin
//			r <= 8'h00;
//			g <= 8'h00;
//			b <= 8'h00;
//		end
//		6: begin
//			r <= 8'h00;
//			g <= 8'h00;
//			b <= 8'h00;
//		7: begin
//			r <= 8'h00;
//			g <= 8'h00;
//			b <= 8'h00;
//		end
//		end
//endmodule
//		