module tb_random_matrix;

    // Parámetros
    reg [3:0] entrada;
    reg [3:0] matriz [7:0][7:0];

    
endmodule
